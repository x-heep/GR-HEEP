../hw/vendor/x-heep/tb/tb_top.sv